`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:53:15 12/10/2022 
// Design Name: 
// Module Name:    ALU_Control_Unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU_Control_Unit(input [2:0]  ALUop , input [5:0]  Function , output reg [3:0] ALUctrl );

	always @(ALUop or Function) begin
			
		if(ALUop == 3'b000) begin
		//------------------------------------------------------------------------------------------------------------
				if(Function == 6'b000000) begin
						assign ALUctrl = 4'b0000;  		//ADD
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000001) begin
						assign ALUctrl = 4'b0001;  		//SUB
					end 
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000010) begin
						assign ALUctrl = 4'b0101;  		//AND
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000011) begin
						assign ALUctrl = 4'b0110;  		//OR
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000100) begin
						assign ALUctrl = 4'b0111;  		//SLT
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000101) begin
						assign ALUctrl = 4'b0011;  		//LSL
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000110) begin
						assign ALUctrl = 4'b0100;  		//LSR
					end
					//------------------------------------------------------------------------------------------------------------
				else if(Function == 6'b000111) begin
						assign ALUctrl = 4'b0010;  		//NOT
					end
					//------------------------------------------------------------------------------------------------------------
			end
			//------------------------------------------------------------------------------------------------------------
		else if(ALUop == 3'b001) begin
				assign ALUctrl = 4'b0001;  				//BEQ SUB
			end
		//------------------------------------------------------------------------------------------------------------
		else if(ALUop == 3'b010) begin
				assign ALUctrl = 4'b0111;  				//SLTI SLT
			end
		//------------------------------------------------------------------------------------------------------------
		else if(ALUop == 3'b011) begin
				assign ALUctrl = 4'b0000;  				//ADDI LW SW  ADD
			end
		//------------------------------------------------------------------------------------------------------------
	end
	//------------------------------------------------------------------------------------------------------------
endmodule
